package fsm_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "trans.sv"
  `include "env_config.sv"

  `include "fsm_seqs.sv"

  `include "driver.sv"
  `include "monitor.sv"
  `include "sequencer.sv"

  `include "agent.sv"

  `include "scoreboard.sv"

  `include "env.sv"

  `include "base_test.sv"

endpackage

