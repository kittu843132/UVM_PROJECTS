package counter_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "trans.sv"
  `include "env_config.sv"

  `include "counter_seqs.sv"

  `include "driver.sv"
  `include "monitor.sv"
  `include "sequencer.sv"

  `include "agent.sv"

  `include "scoreboard.sv"

  `include "env.sv"

  `include "base_test.sv"

endpackage

